library verilog;
use verilog.vl_types.all;
entity alu_test is
end alu_test;
