library verilog;
use verilog.vl_types.all;
entity pc_test is
end pc_test;
