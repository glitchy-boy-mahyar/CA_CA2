library verilog;
use verilog.vl_types.all;
entity shifter_for_jump_test is
end shifter_for_jump_test;
