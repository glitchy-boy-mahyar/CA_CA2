library verilog;
use verilog.vl_types.all;
entity data_mem_test_2 is
end data_mem_test_2;
