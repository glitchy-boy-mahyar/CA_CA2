library verilog;
use verilog.vl_types.all;
entity sign_ext_test is
end sign_ext_test;
