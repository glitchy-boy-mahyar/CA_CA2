library verilog;
use verilog.vl_types.all;
entity data_mem_test is
end data_mem_test;
