library verilog;
use verilog.vl_types.all;
entity inst_mem_test is
end inst_mem_test;
