library verilog;
use verilog.vl_types.all;
entity mux_5bit_test is
end mux_5bit_test;
