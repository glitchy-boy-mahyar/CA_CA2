library verilog;
use verilog.vl_types.all;
entity mux_32bit_test is
end mux_32bit_test;
