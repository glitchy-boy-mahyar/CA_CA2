library verilog;
use verilog.vl_types.all;
entity reg_file_test is
end reg_file_test;
