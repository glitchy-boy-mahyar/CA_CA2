library verilog;
use verilog.vl_types.all;
entity processor_test is
end processor_test;
